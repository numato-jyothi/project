`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:27:18 06/19/2018 
// Design Name: 
// Module Name:    notgate_sim 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created1
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module notgate(a, b);
    input wire a;
    output wire b;
  assign b = !a;


endmodule
